// $Id: $
// File name:   DES_S1.sv
// Created:     4/23/2018
// Author:      Austin Ketterer
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: Sbox 1
module DES_SBOX(input wire [48:1] block, output wire [32:1] out);
   
   wire [3:0] S1[3:0][15:0];
   wire [3:0] S2[3:0][15:0];
   wire [3:0] S3[3:0][15:0];
   wire [3:0] S4[3:0][15:0];
   wire [3:0] S5[3:0][15:0];
   wire [3:0] S6[3:0][15:0];
   wire [3:0] S7[3:0][15:0];
   wire [3:0] S8[3:0][15:0];
   
   assign S1[0][0] = 14;
   assign S1[0][1] = 4;
   assign S1[0][2] = 13;
   assign S1[0][3] = 1;
   assign S1[0][4] = 2;
   assign S1[0][5] = 15;
   assign S1[0][6] = 11;
   assign S1[0][7] = 8;
   assign S1[0][8] = 3;
   assign S1[0][9] = 10;
   assign S1[0][10] = 6;
   assign S1[0][11] = 12;
   assign S1[0][12] = 5;
   assign S1[0][13] = 9;
   assign S1[0][14] = 0;
   assign S1[0][15] = 7;
   assign S1[1][0] = 0;
   assign S1[1][1] = 15;
   assign S1[1][2] = 7;
   assign S1[1][3] = 4;
   assign S1[1][4] = 14;
   assign S1[1][5] = 2;
   assign S1[1][6] = 13;
   assign S1[1][7] = 1;
   assign S1[1][8] = 10;
   assign S1[1][9] = 6;
   assign S1[1][10] = 12;
   assign S1[1][11] = 11;
   assign S1[1][12] = 9;
   assign S1[1][13] = 5;
   assign S1[1][14] = 3;
   assign S1[1][15] = 8;
   assign S1[2][0] = 4;
   assign S1[2][1] = 1;
   assign S1[2][2] = 14;
   assign S1[2][3] = 8;
   assign S1[2][4] = 13;
   assign S1[2][5] = 6;
   assign S1[2][6] = 2;
   assign S1[2][7] = 11;
   assign S1[2][8] = 15;
   assign S1[2][9] = 12;
   assign S1[2][10] = 9;
   assign S1[2][11] = 7;
   assign S1[2][12] = 3;
   assign S1[2][13] = 10;
   assign S1[2][14] = 5;
   assign S1[2][15] = 0;
   assign S1[3][0] = 15;
   assign S1[3][1] = 12;
   assign S1[3][2] = 8;
   assign S1[3][3] = 2;
   assign S1[3][4] = 4;
   assign S1[3][5] = 9;
   assign S1[3][6] = 1;
   assign S1[3][7] = 7;
   assign S1[3][8] = 5;
   assign S1[3][9] = 11;
   assign S1[3][10] = 3;
   assign S1[3][11] = 14;
   assign S1[3][12] = 10;
   assign S1[3][13] = 0;
   assign S1[3][14] = 6;
   assign S1[3][15] = 13;

   assign S2[0][0] = 15;
   assign S2[0][1] = 1;
   assign S2[0][2] = 8;
   assign S2[0][3] = 14;
   assign S2[0][4] = 6;
   assign S2[0][5] = 11;
   assign S2[0][6] = 3;
   assign S2[0][7] = 4;
   assign S2[0][8] = 9;
   assign S2[0][9] = 7;
   assign S2[0][10] = 2;
   assign S2[0][11] = 13;
   assign S2[0][12] = 12;
   assign S2[0][13] = 0;
   assign S2[0][14] = 5;
   assign S2[0][15] = 10;
   assign S2[1][0] = 3;
   assign S2[1][1] = 13;
   assign S2[1][2] = 4;
   assign S2[1][3] = 7;
   assign S2[1][4] = 15;
   assign S2[1][5] = 2;
   assign S2[1][6] = 8;
   assign S2[1][7] = 14;
   assign S2[1][8] = 12;
   assign S2[1][9] = 0;
   assign S2[1][10] = 1;
   assign S2[1][11] = 10;
   assign S2[1][12] = 6;
   assign S2[1][13] = 9;
   assign S2[1][14] = 11;
   assign S2[1][15] = 5;
   assign S2[2][0] = 0;
   assign S2[2][1] = 14;
   assign S2[2][2] = 7;
   assign S2[2][3] = 11;
   assign S2[2][4] = 10;
   assign S2[2][5] = 4;
   assign S2[2][6] = 13;
   assign S2[2][7] = 1;
   assign S2[2][8] = 5;
   assign S2[2][9] = 8;
   assign S2[2][10] = 12;
   assign S2[2][11] = 6;
   assign S2[2][12] = 9;
   assign S2[2][13] = 3;
   assign S2[2][14] = 2;
   assign S2[2][15] = 15;
   assign S2[3][0] = 13;
   assign S2[3][1] = 8;
   assign S2[3][2] = 10;
   assign S2[3][3] = 1;
   assign S2[3][4] = 3;
   assign S2[3][5] = 15;
   assign S2[3][6] = 4;
   assign S2[3][7] = 2;
   assign S2[3][8] = 11;
   assign S2[3][9] = 6;
   assign S2[3][10] = 7;
   assign S2[3][11] = 12;
   assign S2[3][12] = 0;
   assign S2[3][13] = 5;
   assign S2[3][14] = 14;
   assign S2[3][15] = 9;
   assign S3[0][1] = 0;
   assign S3[0][2] = 9;
   assign S3[0][3] = 14;
   assign S3[0][4] = 6;
   assign S3[0][5] = 3;
   assign S3[0][6] = 15;
   assign S3[0][7] = 5;
   assign S3[0][8] = 1;
   assign S3[0][9] = 13;
   assign S3[0][10] = 12;
   assign S3[0][11] = 7;
   assign S3[0][12] = 11;
   assign S3[0][13] = 4;
   assign S3[0][14] = 2;
   assign S3[0][15] = 8;
   assign S3[1][0] = 13;
   assign S3[1][1] = 7;
   assign S3[1][2] = 0;
   assign S3[1][3] = 9;
   assign S3[1][4] = 3;
   assign S3[1][5] = 4;
   assign S3[1][6] = 6;
   assign S3[1][7] = 10;
   assign S3[1][8] = 2;
   assign S3[1][9] = 8;
   assign S3[1][10] = 5;
   assign S3[1][11] = 14;
   assign S3[1][12] = 12;
   assign S3[1][13] = 11;
   assign S3[1][14] = 15;
   assign S3[1][15] = 1;
   assign S3[2][0] = 13;
   assign S3[2][1] = 6;
   assign S3[2][2] = 4;
   assign S3[2][3] = 9;
   assign S3[2][4] = 8;
   assign S3[2][5] = 15;
   assign S3[2][6] = 3;
   assign S3[2][7] = 0;
   assign S3[2][8] = 11;
   assign S3[2][9] = 1;
   assign S3[2][10] = 2;
   assign S3[2][11] = 12;
   assign S3[2][12] = 5;
   assign S3[2][13] = 10;
   assign S3[2][14] = 14;
   assign S3[2][15] = 7;
   assign S3[3][0] = 1;
   assign S3[3][1] = 10;
   assign S3[3][2] = 13;
   assign S3[3][3] = 0;
   assign S3[3][4] = 6;
   assign S3[3][5] = 9;
   assign S3[3][6] = 8;
   assign S3[3][7] = 7;
   assign S3[3][8] = 4;
   assign S3[3][9] = 15;
   assign S3[3][10] = 14;
   assign S3[3][11] = 3;
   assign S3[3][12] = 11;
   assign S3[3][13] = 5;
   assign S3[3][14] = 2;
   assign S3[3][15] = 12;

   assign S4[0][0] = 7;
   assign S4[0][1] = 13;
   assign S4[0][2] = 14;
   assign S4[0][3] = 3;
   assign S4[0][4] = 0;
   assign S4[0][5] = 6;
   assign S4[0][6] = 9;
   assign S4[0][7] = 10;
   assign S4[0][8] = 1;
   assign S4[0][9] = 2;
   assign S4[0][10] = 8;
   assign S4[0][11] = 5;
   assign S4[0][12] = 11;
   assign S4[0][13] = 12;
   assign S4[0][14] = 4;
   assign S4[0][15] = 15;
   assign S4[1][0] = 13;
   assign S4[1][1] = 8;
   assign S4[1][2] = 11;
   assign S4[1][3] = 5;
   assign S4[1][4] = 6;
   assign S4[1][5] = 15;
   assign S4[1][6] = 0;
   assign S4[1][7] = 3;
   assign S4[1][8] = 4;
   assign S4[1][9] = 7;
   assign S4[1][10] = 2;
   assign S4[1][11] = 12;
   assign S4[1][12] = 1;
   assign S4[1][13] = 10;
   assign S4[1][14] = 14;
   assign S4[1][15] = 9;
   assign S4[2][0] = 10;
   assign S4[2][1] = 6;
   assign S4[2][2] = 9;
   assign S4[2][3] = 0;
   assign S4[2][4] = 12;
   assign S4[2][5] = 11;
   assign S4[2][6] = 7;
   assign S4[2][7] = 13;
   assign S4[2][8] = 15;
   assign S4[2][9] = 1;
   assign S4[2][10] = 3;
   assign S4[2][11] = 14;
   assign S4[2][12] = 5;
   assign S4[2][13] = 2;
   assign S4[2][14] = 8;
   assign S4[2][15] = 4;
   assign S4[3][0] = 3;
   assign S4[3][1] = 15;
   assign S4[3][2] = 0;
   assign S4[3][3] = 6;
   assign S4[3][4] = 10;
   assign S4[3][5] = 1;
   assign S4[3][6] = 13;
   assign S4[3][7] = 8;
   assign S4[3][8] = 9;
   assign S4[3][9] = 4;
   assign S4[3][10] = 5;
   assign S4[3][11] = 11;
   assign S4[3][12] = 12;
   assign S4[3][13] = 7;
   assign S4[3][14] = 2;
   assign S4[3][15] = 14;

   assign S5[0][0] = 2;
   assign S5[0][1] = 12;
   assign S5[0][2] = 4;
   assign S5[0][3] = 1;
   assign S5[0][4] = 7;
   assign S5[0][5] = 10;
   assign S5[0][6] = 11;
   assign S5[0][7] = 6;
   assign S5[0][8] = 8;
   assign S5[0][9] = 5;
   assign S5[0][10] = 3;
   assign S5[0][11] = 15;
   assign S5[0][12] = 13;
   assign S5[0][13] = 0;
   assign S5[0][14] = 14;
   assign S5[0][15] = 9;
   assign S5[1][0] = 14;
   assign S5[1][1] = 11;
   assign S5[1][2] = 2;
   assign S5[1][3] = 12;
   assign S5[1][4] = 4;
   assign S5[1][5] = 7;
   assign S5[1][6] = 13;
   assign S5[1][7] = 1;
   assign S5[1][8] = 5;
   assign S5[1][9] = 0;
   assign S5[1][10] = 15;
   assign S5[1][11] = 10;
   assign S5[1][12] = 3;
   assign S5[1][13] = 9;
   assign S5[1][14] = 8;
   assign S5[1][15] = 6;
   assign S5[2][0] = 4;
   assign S5[2][1] = 2;
   assign S5[2][2] = 1;
   assign S5[2][3] = 11;
   assign S5[2][4] = 10;
   assign S5[2][5] = 13;
   assign S5[2][6] = 7;
   assign S5[2][7] = 8;
   assign S5[2][8] = 15;
   assign S5[2][9] = 9;
   assign S5[2][10] = 12;
   assign S5[2][11] = 5;
   assign S5[2][12] = 6;
   assign S5[2][13] = 3;
   assign S5[2][14] = 0;
   assign S5[2][15] = 14;
   assign S5[3][0] = 11;
   assign S5[3][1] = 8;
   assign S5[3][2] = 12;
   assign S5[3][3] = 7;
   assign S5[3][4] = 1;
   assign S5[3][5] = 14;
   assign S5[3][6] = 2;
   assign S5[3][7] = 13;
   assign S5[3][8] = 6;
   assign S5[3][9] = 15;
   assign S5[3][10] = 0;
   assign S5[3][11] = 9;
   assign S5[3][12] = 10;
   assign S5[3][13] = 4;
   assign S5[3][14] = 5;
   assign S5[3][15] = 3;

   assign S6[0][0] = 12;
   assign S6[0][1] = 1;
   assign S6[0][2] = 10;
   assign S6[0][3] = 15;
   assign S6[0][4] = 9;
   assign S6[0][5] = 2;
   assign S6[0][6] = 6;
   assign S6[0][7] = 8;
   assign S6[0][8] = 0;
   assign S6[0][9] = 13;
   assign S6[0][10] = 3;
   assign S6[0][11] = 4;
   assign S6[0][12] = 14;
   assign S6[0][13] = 7;
   assign S6[0][14] = 5;
   assign S6[0][15] = 11;
   assign S6[1][0] = 10;
   assign S6[1][1] = 15;
   assign S6[1][2] = 4;
   assign S6[1][3] = 2;
   assign S6[1][4] = 7;
   assign S6[1][5] = 12;
   assign S6[1][6] = 9;
   assign S6[1][7] = 5;
   assign S6[1][8] = 6;
   assign S6[1][9] = 1;
   assign S6[1][10] = 13;
   assign S6[1][11] = 14;
   assign S6[1][12] = 0;
   assign S6[1][13] = 11;
   assign S6[1][14] = 3;
   assign S6[1][15] = 8;
   assign S6[2][0] = 9;
   assign S6[2][1] = 14;
   assign S6[2][2] = 15;
   assign S6[2][3] = 5;
   assign S6[2][4] = 2;
   assign S6[2][5] = 8;
   assign S6[2][6] = 12;
   assign S6[2][7] = 3;
   assign S6[2][8] = 7;
   assign S6[2][9] = 0;
   assign S6[2][10] = 4;
   assign S6[2][11] = 10;
   assign S6[2][12] = 1;
   assign S6[2][13] = 13;
   assign S6[2][14] = 11;
   assign S6[2][15] = 6;
   assign S6[3][0] = 4;
   assign S6[3][1] = 3;
   assign S6[3][2] = 2;
   assign S6[3][3] = 12;
   assign S6[3][4] = 9;
   assign S6[3][5] = 5;
   assign S6[3][6] = 15;
   assign S6[3][7] = 10;
   assign S6[3][8] = 11;
   assign S6[3][9] = 14;
   assign S6[3][10] = 1;
   assign S6[3][11] = 7;
   assign S6[3][12] = 6;
   assign S6[3][13] = 0;
   assign S6[3][14] = 8;
   assign S6[3][15] = 13;

   assign S7[0][0] = 4;
   assign S7[0][1] = 11;
   assign S7[0][2] = 2;
   assign S7[0][3] = 14;
   assign S7[0][4] = 15;
   assign S7[0][5] = 0;
   assign S7[0][6] = 8;
   assign S7[0][7] = 13;
   assign S7[0][8] = 3;
   assign S7[0][9] = 12;
   assign S7[0][10] = 9;
   assign S7[0][11] = 7;
   assign S7[0][12] = 5;
   assign S7[0][13] = 10;
   assign S7[0][14] = 6;
   assign S7[0][15] = 1;
   assign S7[1][0] = 13;
   assign S7[1][1] = 0;
   assign S7[1][2] = 11;
   assign S7[1][3] = 7;
   assign S7[1][4] = 4;
   assign S7[1][5] = 9;
   assign S7[1][6] = 1;
   assign S7[1][7] = 10;
   assign S7[1][8] = 14;
   assign S7[1][9] = 3;
   assign S7[1][10] = 5;
   assign S7[1][11] = 12;
   assign S7[1][12] = 2;
   assign S7[1][13] = 15;
   assign S7[1][14] = 8;
   assign S7[1][15] = 6;
   assign S7[2][0] = 1;
   assign S7[2][1] = 4;
   assign S7[2][2] = 11;
   assign S7[2][3] = 13;
   assign S7[2][4] = 12;
   assign S7[2][5] = 3;
   assign S7[2][6] = 7;
   assign S7[2][7] = 14;
   assign S7[2][8] = 10;
   assign S7[2][9] = 15;
   assign S7[2][10] = 6;
   assign S7[2][11] = 8;
   assign S7[2][12] = 0;
   assign S7[2][13] = 5;
   assign S7[2][14] = 9;
   assign S7[2][15] = 2;
   assign S7[3][0] = 6;
   assign S7[3][1] = 11;
   assign S7[3][2] = 13;
   assign S7[3][3] = 8;
   assign S7[3][4] = 1;
   assign S7[3][5] = 4;
   assign S7[3][6] = 10;
   assign S7[3][7] = 7;
   assign S7[3][8] = 9;
   assign S7[3][9] = 5;
   assign S7[3][10] = 0;
   assign S7[3][11] = 15;
   assign S7[3][12] = 14;
   assign S7[3][13] = 2;
   assign S7[3][14] = 3;
   assign S7[3][15] = 12;

   assign S8[0][0] = 13;
   assign S8[0][1] = 2;
   assign S8[0][2] = 8;
   assign S8[0][3] = 4;
   assign S8[0][4] = 6;
   assign S8[0][5] = 15;
   assign S8[0][6] = 11;
   assign S8[0][7] = 1;
   assign S8[0][8] = 10;
   assign S8[0][9] = 9;
   assign S8[0][10] = 3;
   assign S8[0][11] = 14;
   assign S8[0][12] = 5;
   assign S8[0][13] = 0;
   assign S8[0][14] = 12;
   assign S8[0][15] = 7;
   assign S8[1][0] = 1;
   assign S8[1][1] = 15;
   assign S8[1][2] = 13;
   assign S8[1][3] = 8;
   assign S8[1][4] = 10;
   assign S8[1][5] = 3;
   assign S8[1][6] = 7;
   assign S8[1][7] = 4;
   assign S8[1][8] = 12;
   assign S8[1][9] = 5;
   assign S8[1][10] = 6;
   assign S8[1][11] = 11;
   assign S8[1][12] = 0;
   assign S8[1][13] = 14;
   assign S8[1][14] = 9;
   assign S8[1][15] = 2;
   assign S8[2][0] = 7;
   assign S8[2][1] = 11;
   assign S8[2][2] = 4;
   assign S8[2][3] = 1;
   assign S8[2][4] = 9;
   assign S8[2][5] = 12;
   assign S8[2][6] = 14;
   assign S8[2][7] = 2;
   assign S8[2][8] = 0;
   assign S8[2][9] = 6;
   assign S8[2][10] = 10;
   assign S8[2][11] = 13;
   assign S8[2][12] = 15;
   assign S8[2][13] = 3;
   assign S8[2][14] = 5;
   assign S8[2][15] = 8;
   assign S8[3][0] = 2;
   assign S8[3][1] = 1;
   assign S8[3][2] = 14;
   assign S8[3][3] = 7;
   assign S8[3][4] = 4;
   assign S8[3][5] = 10;
   assign S8[3][6] = 8;
   assign S8[3][7] = 13;
   assign S8[3][8] = 15;
   assign S8[3][9] = 12;
   assign S8[3][10] = 9;
   assign S8[3][11] = 0;
   assign S8[3][12] = 3;
   assign S8[3][13] = 5;
   assign S8[3][14] = 6;
   assign S8[3][15] = 11;

   assign out[32:29] = S1[{block[48], block[43]}][block[47:44]];
   assign out[28:25] = S2[{block[42], block[37]}][block[41:38]];
   assign out[24:21] = S3[{block[36], block[31]}][block[35:32]];
   assign out[20:17] = S4[{block[30], block[25]}][block[29:26]];
   assign out[16:13] = S5[{block[24], block[19]}][block[23:20]];
   assign out[12:9] = S6[{block[18], block[13]}][block[17:14]];
   assign out[8:5]  = S7[{block[12], block[7]}][block[11:8]];
   assign out[4:1]   = S8[{block[6], block[1]}][block[5:2]];
endmodule // DES_S1

