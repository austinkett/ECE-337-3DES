// $Id: $
// File name:   tb_DES_flex_counter.sv
// Created:     4/23/2018
// Author:      Austin Ketterer
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: tb for flex
